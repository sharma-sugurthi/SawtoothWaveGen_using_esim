* C:\Users\PC\eSim-Workspace\Triangular\Triangular.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 2/9/2025 6:02:41 PM

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
X1  ? GND Net-_R1-Pad1_ Net-_X1-Pad4_ ? out1 Net-_X1-Pad7_ ? lm_741		
X2  ? Net-_C1-Pad2_ GND Net-_X1-Pad4_ ? out2 Net-_X1-Pad7_ ? lm_741		
v1  GND Net-_X1-Pad4_ 14V		
v2  Net-_X1-Pad7_ GND 14V		
R2  Net-_R1-Pad1_ out1 1k		
R3  out1 Net-_C1-Pad2_ 10k		
R1  Net-_R1-Pad1_ out2 180		
U2  out2 plot_v1		
U1  out1 plot_v1		
C1  out2 Net-_C1-Pad2_ 47n		

.end
