* C:\Users\PC\eSim-Workspace\Sawtooth\Sawtooth.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 2/10/2025 11:01:08 AM

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
X1  ? GND Net-_R1-Pad2_ Net-_X1-Pad4_ ? out1 Net-_X1-Pad7_ ? lm_741		
X2  ? Net-_C1-Pad2_ GND Net-_X1-Pad4_ ? out2 Net-_X1-Pad7_ ? lm_741		
R3  Net-_D2-Pad2_ Net-_C1-Pad2_ 5k		
R2  Net-_R1-Pad2_ out2 40k		
R1  out1 Net-_R1-Pad2_ 100k		
R4  Net-_D1-Pad1_ Net-_C1-Pad2_ 40k		
v2  GND Net-_X1-Pad4_ 15V		
v1  Net-_X1-Pad7_ GND 15V		
D2  out1 Net-_D2-Pad2_ eSim_Diode		
D1  Net-_D1-Pad1_ out1 eSim_Diode		
C1  out2 Net-_C1-Pad2_ 500nF		
U2  out2 plot_v1		
U1  out1 plot_v1		

.end
